interface intf ();
    // STEP 1: define your interface signals here
    logic clk;
    logic reset_n;
    logic d_in;
    logic q_out;
endinterface : intf
