interface intf ();
    // STEP 1: define your interface signals here
endinterface : intf
