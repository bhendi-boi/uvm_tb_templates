interface intf ();
	// input ports
	logic clk;
	logic reset_n;
	logic d_in;

	// output ports
	logic q_out;
endinterface : intf
